0
0 0 0 0 0 g c 4 1 34 1
0 0 0 0 0 g c 6 1 23 1
0 0 0 0 0 g c 8 1 32 1
0 0 0 0 0 g c 45 1 36 1
1 10 4 8 0 9 5 7 3 9 4 8 0 6 4 10 1 12 3 6 3 5 2 2 0 3 2 11 0 5 2 3 1 4 2 11 1 4 
